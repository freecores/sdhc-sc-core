//
// file: SDCommandArg.sv
// author: Rainer Kastl
//
// 
//
 
`ifndef SDCOMMANDARG
`define SDCOMMANDARG

`define cSDArgWith 32
typedef logic[`cSDArgWith-1:0] SDCommandArg;

`endif
