`ifndef RAMACTION_SV
`define RAMACTION_SV

class RamAction;

endclass

typedef mailbox #(RamAction) RamActionMb;

`endif

