`ifndef EXPECTEDRESULT_SV
`define EXPECTEDRESULT_SV

class ExpectedResult;
endclass

typedef mailbox #(ExpectedResult) ExpectedResultMb;

`endif
