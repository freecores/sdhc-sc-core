`ifndef SDCORETRANSACTIONBFM_SV
`define SDCORETRANSACTIONBFM_SV

class SdCoreTransactionBFM;

endclass

`endif
