`ifndef SDCORETRANSFERFUNCTION_SV
`define SDCORETRANSFERFUNCTION_SV

`include "SdCoreTransaction.sv";

class SdCoreTransferFunction;
	SdCoreTransSeqMb TransInMb;

endclass

`endif
