
`ifndef WBTRANSACTION_SV
`define WBTRANSACTION_SV

class WbTransaction;
endclass

typedef mailbox #(WbTransaction) WbTransMb;

`endif

