`ifndef SDCORECHECKER_SV
`define SDCORECHECKER_SV

class SdCoreChecker;

endclass

`endif
